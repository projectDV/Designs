/********************************************************************************************
Copyright 2019 - Maven Silicon Softech Pvt Ltd. 
 
All Rights Reserved.

This source code is an unpublished work belongs to Maven Silicon Softech Pvt Ltd.

It is not to be shared with or used by any third parties who have not enrolled for our paid training 

courses or received any written authorization from Maven Silicon.


Webpage:  www.maven-silicon.com

Filename:	  mux4_1.v   

Description:      4:1 Mux Design

Author Name:       Susmita

Version: 1.0
*********************************************************************************************/
 
module mux4_1(input a,b,c,d,
              s1,s0,
              output y);


// Step 1. Declare the internal wires
 

// Step 2. Instantiate the 2:1 Mux and map the ports


endmodule
  

module mux4_1(input a,b,c,d,
              s1,s0,
              output y);

endmodule
  
